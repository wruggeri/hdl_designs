/*
File name:      apb_parameters.svh
Author:         Walter Ruggeri
Description:    parameters to configure an APB slave and its test environment

28/08/2022      Initial release
*/


localparam N_BIT_DATA = 32;
localparam N_BIT_ADDRESS = 8;
localparam DELAY_NS = 27;
localparam CLOCK_PERIOD_NS = 10;